module DDS_FIR(
    input wire clk,
   );
endmodule